module order_quantity #
(
   input logic i_clk,
   input logic 
)
(
    
);
    
   
endmodule
