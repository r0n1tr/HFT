// This file is public domain, it can be freely copied without restrictions.
// SPDX-License-Identifier: CC0-1.0


module my_design
(
    input logic clk,
    output logic my_signal_1,
    output logic my_signal_2
);


  assign my_signal_1 = 1'bx;
  assign my_signal_2 = 0;


endmodule
